--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   03:44:05 03/10/2022
-- Design Name:   
-- Module Name:   G:/xlinx_projects/computer_arch/LAB1/sipo_test.vhd
-- Project Name:  LAB1
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: sipo
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY sipo_test IS
END sipo_test;
 
ARCHITECTURE behavior OF sipo_test IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT sipo
    PORT(
         clk : IN  std_logic;
         A : IN  std_logic;
         SHIFTA : IN  std_logic;
         A_out : OUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal A : std_logic := '0';
   signal SHIFTA : std_logic := '0';

 	--Outputs
   signal A_out : std_logic_vector(3 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: sipo PORT MAP (
          clk => clk,
          A => A,
          SHIFTA => SHIFTA,
          A_out => A_out
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 10 ns;	
		A<='0';
		SHIFTA<='1';
		wait for 10 ns;
		A<='1';
		SHIFTA<='1';
		wait for 10 ns;
		A<='1';
		SHIFTA<='1';
		wait for 10 ns;
		A<='0';
		SHIFTA<='1';
		wait for 10 ns;
		A<='1';
		SHIFTA<='1';
		wait for 10 ns;
		A<='1';
		SHIFTA<='1';
		wait for 10 ns;
		A<='0';
		SHIFTA<='1';
		wait for 10 ns;
		A<='0';
      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
